vpalladi@outatime.cern.ch.19264:1548249750